//TODO: MAKE THE TOP MODULE
